`timescale 1ns / 1ps
`include "params.vh"

module element_wise #
(

)
(

);

endmodule  // element_wise