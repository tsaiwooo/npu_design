// 目前的問題是axi_stream_output的tvalid跟start_output不一樣導致addr錯誤, 取到錯的data, 還有存入sram的data有幾個也是錯的需要去debug
`timescale 1ns / 1ps
`include "params.vh"

module npu #
(
    parameter MAX_MACS = 64,
    parameter ADDR_WIDTH = 13,
    parameter C_AXIS_TDATA_WIDTH = 8,
    parameter C_AXIS_MDATA_WIDTH = 8,
    parameter MAX_CHANNELS = 64,
    parameter NUM_CHANNELS_WIDTH = $clog2(MAX_CHANNELS+1),
    parameter QUANT_WIDTH = 32
)
(
    /* AXI slave interface (input to the FIFO) */
    input  wire                   s00_axis_aclk,
    input  wire                   s00_axis_aresetn,
    input  wire signed [C_AXIS_TDATA_WIDTH-1:0]  s00_axis_tdata,
    input  wire [(C_AXIS_TDATA_WIDTH/8)-1 : 0]   s00_axis_tstrb,
    input  wire                   s00_axis_tvalid,
    output wire                   s00_axis_tready,
    input  wire                   s00_axis_tlast,
    input  wire [2*ADDR_WIDTH + NUM_CHANNELS_WIDTH-1:0] s00_axis_tuser,  

    /* AXI master interface (output of the FIFO) */
    input  wire                   m00_axis_aclk,
    input  wire                   m00_axis_aresetn,
    output wire signed [4*C_AXIS_MDATA_WIDTH-1:0]  m00_axis_tdata,
    output wire [(2*C_AXIS_MDATA_WIDTH/8)-1 : 0]   m00_axis_tstrb, 
    output wire                   m00_axis_tvalid,
    input  wire                   m00_axis_tready,
    output wire                   m00_axis_tlast,
    output wire [NUM_CHANNELS_WIDTH-1:0]           m00_axis_tuser, 

    // requant signals
    input wire [31:0]            quantized_multiplier,
    input wire signed  [31:0]     shift


);

    reg [2:0] state = IDLE, next_state;
    reg start_output = 1'b0;
    reg GEMM_en = 1'b0;
    reg ELEMENT_en = 1'b0;

    // axi_stream_input signals
    wire                    write_enable;
    wire [ADDR_WIDTH-1:0]   write_address;
    wire signed [C_AXIS_TDATA_WIDTH-1:0] write_data;
    wire [2:0]              data_type;
    wire                    data_ready;
    wire [ADDR_WIDTH-1:0]   img_row;
    wire [ADDR_WIDTH-1:0]   img_col;
    wire [ADDR_WIDTH-1:0]   ker_row;
    wire [ADDR_WIDTH-1:0]   ker_col;
    wire [NUM_CHANNELS_WIDTH-1:0] num_channels;


    // axi_stream_output signals
    wire                   sram_out_en;
    wire [MAX_ADDR_WIDTH-1:0]  sram_out_addr;

    // convolution signals
    wire signed [C_AXIS_MDATA_WIDTH - 1 : 0] mac_out;
    wire mac_valid_out;

    // output index control
    wire [MAX_ADDR_WIDTH-1:0] idx1_out;

    // output size
    wire [ADDR_WIDTH-1:0] out_row, out_col;
    assign out_row = img_row - ker_row + 1;
    assign out_col = img_col - ker_col + 1;


    // GEMM convolution index
    wire [ADDR_WIDTH-1:0] conv_row;
    wire [ADDR_WIDTH-1:0] conv_col;
    wire [ADDR_WIDTH-1:0] for_conv_row;
    wire [ADDR_WIDTH-1:0] for_conv_col;
    wire [ADDR_WIDTH-1:0] weight_idx;


    // SRAM OUTPUT DATA
    wire signed [SRAM_WIDTH_O-1:0] gemm0_data_out;
    wire signed [SRAM_WIDTH_O-1:0] gemm1_data_out;
    wire signed [SRAM_WIDTH_O-1:0] elem_data_out;
    wire signed [SRAM_WIDTH_O-1:0] sram_data_out;

    // requant signals
    wire requant_valid_o;

    // control FSM
    always @(*) begin
        next_state = state;
        case (state)
            IDLE: begin
                if (data_ready && data_type == GEMM0_SRAM_IDX)
                    next_state = LOAD_IMG;
            end
            LOAD_IMG: begin
                if (data_ready && data_type == GEMM1_SRAM_IDX)
                    next_state = LOAD_KER;
            end
            LOAD_KER: begin
                // assum that the data is ready
                if (!data_ready)
                    next_state = COMPUTE_CONV0;
            end
            COMPUTE_CONV0: begin
                // if (conv_row >= out_row - 1 && conv_col >= out_col - 1 && for_conv_row == ker_row) begin
                //     next_state = WAIT_LAST;
                // end else if (for_conv_row == ker_row ) begin
                //     next_state = COMPUTE_CONV1;
                // end else begin
                //     next_state = COMPUTE_CONV0;
                // end
                next_state = (start_output)? WRITE_OUTPUT : COMPUTE_CONV0;
            end
            // COMPUTE_CONV1: begin
            //     next_state = COMPUTE_CONV0;
            // end
            // WAIT_LAST: begin
            //     if (mac_valid_out)
            //         next_state = WRITE_OUTPUT;
            // end
            WRITE_OUTPUT: begin
                if (sram_out_addr >= out_row * out_col)begin
                    next_state = IDLE;
                end 
            end
            default: next_state = IDLE;
        endcase
    end

    always @(posedge s00_axis_aclk) begin
        if (!s00_axis_aresetn)begin
            state <= IDLE;
        end else begin
            state <= next_state;
        end
    end
    
    // control GEMM_en
    always @(posedge s00_axis_aclk)begin
        if(!s00_axis_aresetn)begin
            GEMM_en <= 1'b0;
        end else if(conv_row == out_row)begin
            GEMM_en <= 1'b0;
        end else if(state == COMPUTE_CONV0)begin
            GEMM_en <= 1'b1;
        end else if(idx1_out == (out_col * out_row -1))begin
            GEMM_en <= 1'b0;
        end
    end

    // control start_output
    always @(posedge s00_axis_aclk)begin
        if(!s00_axis_aresetn)begin
            start_output <= 1'b0;
        end else if(idx1_out == (out_col * out_row -1) && state == COMPUTE_CONV0)begin
            start_output <= 1'b1;
        end
    end

    GEMM #
    (
        .MAX_MACS(MAX_MACS),
        .ADDR_WIDTH(ADDR_WIDTH),
        .DATA_WIDTH(C_AXIS_TDATA_WIDTH)
    )
    GEMM_inst
    (
        .clk(s00_axis_aclk),
        .rst(s00_axis_aresetn),
        // convolution signals
        .convolution_en(GEMM_en),
        // input metadata
        .img_row(img_row),
        .img_col(img_col),
        .ker_row(ker_row),
        .ker_col(ker_col),
        // img and kernel data
        .data_in(gemm0_data_out),
        .weight_in(gemm1_data_out),
        // output signal control
        .mac_valid_out(mac_valid_out),
        .mac_out(mac_out),
        // output metadata
        .conv_row(conv_row),
        .conv_col(conv_col),
        .for_conv_row(for_conv_row),
        .for_conv_col(for_conv_col),
        .weight_idx_o(weight_idx),
        // quantized multiplier and shift given by testbench temporarily
        .quantized_multiplier(quantized_multiplier),
        .shift(shift),
        .requant_valid_o(requant_valid_o),
        .idx1_out(idx1_out)
    );


    axi_stream_input #
    (
        .ADDR_WIDTH(ADDR_WIDTH),
        .DATA_WIDTH(C_AXIS_TDATA_WIDTH),
        .NUM_CHANNELS_WIDTH(NUM_CHANNELS_WIDTH)
    )
    axi_stream_input_inst
    (
        .s_axis_aclk(s00_axis_aclk),
        .s_axis_aresetn(s00_axis_aresetn),
        .s_axis_tdata(s00_axis_tdata),
        .s_axis_tstrb(s00_axis_tstrb),
        .s_axis_tvalid(s00_axis_tvalid),
        .s_axis_tready(s00_axis_tready),
        .s_axis_tlast(s00_axis_tlast),
        .s_axis_tuser(s00_axis_tuser),
        .write_enable(write_enable),
        .write_address(write_address),
        .write_data(write_data),
        .data_type(data_type),
        .data_ready(data_ready),
        .img_row(img_row),
        .img_col(img_col),
        .ker_row(ker_row),
        .ker_col(ker_col),
        .num_channels(num_channels)
    );


    axi_stream_output #
    (
        .ADDR_WIDTH(ADDR_WIDTH),
        .DATA_WIDTH(C_AXIS_MDATA_WIDTH),
        .NUM_CHANNELS_WIDTH(NUM_CHANNELS_WIDTH)
    )
    axi_stream_output_inst
    (
        .m_axis_aclk(m00_axis_aclk),
        .m_axis_aresetn(m00_axis_aresetn),
        .m_axis_tdata(m00_axis_tdata),
        // .m_axis_tstrb(m00_axis_tstrb),
        .m_axis_tvalid(m00_axis_tvalid),
        .m_axis_tready(m00_axis_tready),
        .m_axis_tlast(m00_axis_tlast),
        .m_axis_tuser(m00_axis_tuser),
        // SRAM interface
        .sram_out_en(sram_out_en),
        .sram_out_addr(sram_out_addr),
        .sram_out_data_out(sram_data_out),
        // control signals
        .start_output(state == WRITE_OUTPUT),
        .out_size(out_row * out_col)
    );

    sram_controller sram_controller_inst
    (
        .clk(s00_axis_aclk),
        .rst(s00_axis_aresetn),
        // GEMM1 port
        .gemm1_addr((conv_row + for_conv_row) * img_col + conv_col + for_conv_col),
        .gemm1_data_in(),
        .gemm1_en(state == COMPUTE_CONV0),
        .gemm1_we(1'b0),
        .gemm1_idx(GEMM0_SRAM_IDX),
        .gemm1_data_out(gemm0_data_out),
        // GEMM2 port
        .gemm2_addr(weight_idx),
        .gemm2_data_in(),
        .gemm2_en(state == COMPUTE_CONV0),
        .gemm2_we(1'b0),
        .gemm2_idx(GEMM1_SRAM_IDX),
        .gemm2_data_out(gemm1_data_out),
        // ELEM port
        .elem_addr(idx1_out),
        .elem_data_in(mac_out),
        // .elem_en(mac_valid_out),
        // .elem_we(mac_valid_out),
        .elem_en(requant_valid_o),
        .elem_we(requant_valid_o),
        .elem_idx(ELEM0_SRAM_IDX),
        .elem_data_out(elem_data_out),
        // axi4 input port
        .write_address(write_address),
        .write_data(write_data),
        .axi_idx(data_type),
        .write_enable(write_enable),
        // axi4 output port
        .sram_out_en(sram_out_en),
        .sram_out_idx(ELEM0_SRAM_IDX),
        .sram_out_addr(sram_out_addr),
        .sram_out_data(sram_data_out)
    );

endmodule
